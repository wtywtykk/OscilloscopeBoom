Package ScanParam Is
	Constant VGADimensionBits:INTEGER:=13;
	Constant LineMinScanTime:INTEGER:=4801;
	Constant ScanLeft:INTEGER:=200;
	Constant ScanTop:INTEGER:=200;
	Constant ScanWidth:INTEGER:=400;
	Constant ScanHeight:INTEGER:=300;
	Constant MemAddrBits:INTEGER:=17;
	Constant PixelBits:INTEGER:=4;
	Constant ScanPixelBits:INTEGER:=13;
End ScanParam;
